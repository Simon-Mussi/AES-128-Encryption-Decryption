// Inverse SBox module for decryption.
module INV_SBOX(
    input clk,
    input [7:0] IN_DATA,
    output [7:0] OUT_DATA
  );
  
    reg [7:0] OUT_REG;
    // Perform substitution based on the predefined inverse AES SBox table.
    always @(posedge clk) begin
      case (IN_DATA)
        8'h00: OUT_REG <= 8'h52;
        8'h01: OUT_REG <= 8'h09;
        8'h02: OUT_REG <= 8'h6a;
        8'h03: OUT_REG <= 8'hd5;
        8'h04: OUT_REG <= 8'h30;
        8'h05: OUT_REG <= 8'h36;
        8'h06: OUT_REG <= 8'ha5;
        8'h07: OUT_REG <= 8'h38;
        8'h08: OUT_REG <= 8'hbf;
        8'h09: OUT_REG <= 8'h40;
        8'h0a: OUT_REG <= 8'ha3;
        8'h0b: OUT_REG <= 8'h9e;
        8'h0c: OUT_REG <= 8'h81;
        8'h0d: OUT_REG <= 8'hf3;
        8'h0e: OUT_REG <= 8'hd7;
        8'h0f: OUT_REG <= 8'hfb;
        8'h10: OUT_REG <= 8'h7c;
        8'h11: OUT_REG <= 8'he3;
        8'h12: OUT_REG <= 8'h39;
        8'h13: OUT_REG <= 8'h82;
        8'h14: OUT_REG <= 8'h9b;
        8'h15: OUT_REG <= 8'h2f;
        8'h16: OUT_REG <= 8'hff;
        8'h17: OUT_REG <= 8'h87;
        8'h18: OUT_REG <= 8'h34;
        8'h19: OUT_REG <= 8'h8e;
        8'h1a: OUT_REG <= 8'h43;
        8'h1b: OUT_REG <= 8'h44;
        8'h1c: OUT_REG <= 8'hc4;
        8'h1d: OUT_REG <= 8'hde;
        8'h1e: OUT_REG <= 8'he9;
        8'h1f: OUT_REG <= 8'hcb;
        8'h20: OUT_REG <= 8'h54;
        8'h21: OUT_REG <= 8'h7b;
        8'h22: OUT_REG <= 8'h94;
        8'h23: OUT_REG <= 8'h32;
        8'h24: OUT_REG <= 8'ha6;
        8'h25: OUT_REG <= 8'hc2;
        8'h26: OUT_REG <= 8'h23;
        8'h27: OUT_REG <= 8'h3d;
        8'h28: OUT_REG <= 8'hee;
        8'h29: OUT_REG <= 8'h4c;
        8'h2a: OUT_REG <= 8'h95;
        8'h2b: OUT_REG <= 8'h0b;
        8'h2c: OUT_REG <= 8'h42;
        8'h2d: OUT_REG <= 8'hfa;
        8'h2e: OUT_REG <= 8'hc3;
        8'h2f: OUT_REG <= 8'h4e;
        8'h30: OUT_REG <= 8'h08;
        8'h31: OUT_REG <= 8'h2e;
        8'h32: OUT_REG <= 8'ha1;
        8'h33: OUT_REG <= 8'h66;
        8'h34: OUT_REG <= 8'h28;
        8'h35: OUT_REG <= 8'hd9;
        8'h36: OUT_REG <= 8'h24;
        8'h37: OUT_REG <= 8'hb2;
        8'h38: OUT_REG <= 8'h76;
        8'h39: OUT_REG <= 8'h5b;
        8'h3a: OUT_REG <= 8'ha2;
        8'h3b: OUT_REG <= 8'h49;
        8'h3c: OUT_REG <= 8'h6d;
        8'h3d: OUT_REG <= 8'h8b;
        8'h3e: OUT_REG <= 8'hd1;
        8'h3f: OUT_REG <= 8'h25;
        8'h40: OUT_REG <= 8'h72;
        8'h41: OUT_REG <= 8'hf8;
        8'h42: OUT_REG <= 8'hf6;
        8'h43: OUT_REG <= 8'h64;
        8'h44: OUT_REG <= 8'h86;
        8'h45: OUT_REG <= 8'h68;
        8'h46: OUT_REG <= 8'h98;
        8'h47: OUT_REG <= 8'h16;
        8'h48: OUT_REG <= 8'hd4;
        8'h49: OUT_REG <= 8'ha4;
        8'h4a: OUT_REG <= 8'h5c;
        8'h4b: OUT_REG <= 8'hcc;
        8'h4c: OUT_REG <= 8'h5d;
        8'h4d: OUT_REG <= 8'h65;
        8'h4e: OUT_REG <= 8'hb6;
        8'h4f: OUT_REG <= 8'h92;
        8'h50: OUT_REG <= 8'h6c;
        8'h51: OUT_REG <= 8'h70;
        8'h52: OUT_REG <= 8'h48;
        8'h53: OUT_REG <= 8'h50;
        8'h54: OUT_REG <= 8'hfd;
        8'h55: OUT_REG <= 8'hed;
        8'h56: OUT_REG <= 8'hb9;
        8'h57: OUT_REG <= 8'hda;
        8'h58: OUT_REG <= 8'h5e;
        8'h59: OUT_REG <= 8'h15;
        8'h5a: OUT_REG <= 8'h46;
        8'h5b: OUT_REG <= 8'h57;
        8'h5c: OUT_REG <= 8'ha7;
        8'h5d: OUT_REG <= 8'h8d;
        8'h5e: OUT_REG <= 8'h9d;
        8'h5f: OUT_REG <= 8'h84;
        8'h60: OUT_REG <= 8'h90;
        8'h61: OUT_REG <= 8'hd8;
        8'h62: OUT_REG <= 8'hab;
        8'h63: OUT_REG <= 8'h00;
        8'h64: OUT_REG <= 8'h8c;
        8'h65: OUT_REG <= 8'hbc;
        8'h66: OUT_REG <= 8'hd3;
        8'h67: OUT_REG <= 8'h0a;
        8'h68: OUT_REG <= 8'hf7;
        8'h69: OUT_REG <= 8'he4;
        8'h6a: OUT_REG <= 8'h58;
        8'h6b: OUT_REG <= 8'h05;
        8'h6c: OUT_REG <= 8'hb8;
        8'h6d: OUT_REG <= 8'hb3;
        8'h6e: OUT_REG <= 8'h45;
        8'h6f: OUT_REG <= 8'h06;
        8'h70: OUT_REG <= 8'hd0;
        8'h71: OUT_REG <= 8'h2c;
        8'h72: OUT_REG <= 8'h1e;
        8'h73: OUT_REG <= 8'h8f;
        8'h74: OUT_REG <= 8'hca;
        8'h75: OUT_REG <= 8'h3f;
        8'h76: OUT_REG <= 8'h0f;
        8'h77: OUT_REG <= 8'h02;
        8'h78: OUT_REG <= 8'hc1;
        8'h79: OUT_REG <= 8'haf;
        8'h7a: OUT_REG <= 8'hbd;
        8'h7b: OUT_REG <= 8'h03;
        8'h7c: OUT_REG <= 8'h01;
        8'h7d: OUT_REG <= 8'h13;
        8'h7e: OUT_REG <= 8'h8a;
        8'h7f: OUT_REG <= 8'h6b;
        8'h80: OUT_REG <= 8'h3a;
        8'h81: OUT_REG <= 8'h91;
        8'h82: OUT_REG <= 8'h11;
        8'h83: OUT_REG <= 8'h41;
        8'h84: OUT_REG <= 8'h4f;
        8'h85: OUT_REG <= 8'h67;
        8'h86: OUT_REG <= 8'hdc;
        8'h87: OUT_REG <= 8'hea;
        8'h88: OUT_REG <= 8'h97;
        8'h89: OUT_REG <= 8'hf2;
        8'h8a: OUT_REG <= 8'hcf;
        8'h8b: OUT_REG <= 8'hce;
        8'h8c: OUT_REG <= 8'hf0;
        8'h8d: OUT_REG <= 8'hb4;
        8'h8e: OUT_REG <= 8'he6;
        8'h8f: OUT_REG <= 8'h73;
        8'h90: OUT_REG <= 8'h96;
        8'h91: OUT_REG <= 8'hac;
        8'h92: OUT_REG <= 8'h74;
        8'h93: OUT_REG <= 8'h22;
        8'h94: OUT_REG <= 8'he7;
        8'h95: OUT_REG <= 8'had;
        8'h96: OUT_REG <= 8'h35;
        8'h97: OUT_REG <= 8'h85;
        8'h98: OUT_REG <= 8'he2;
        8'h99: OUT_REG <= 8'hf9;
        8'h9a: OUT_REG <= 8'h37;
        8'h9b: OUT_REG <= 8'he8;
        8'h9c: OUT_REG <= 8'h1c;
        8'h9d: OUT_REG <= 8'h75;
        8'h9e: OUT_REG <= 8'hdf;
        8'h9f: OUT_REG <= 8'h6e;
        8'ha0: OUT_REG <= 8'h47;
        8'ha1: OUT_REG <= 8'hf1;
        8'ha2: OUT_REG <= 8'h1a;
        8'ha3: OUT_REG <= 8'h71;
        8'ha4: OUT_REG <= 8'h1d;
        8'ha5: OUT_REG <= 8'h29;
        8'ha6: OUT_REG <= 8'hc5;
        8'ha7: OUT_REG <= 8'h89;
        8'ha8: OUT_REG <= 8'h6f;
        8'ha9: OUT_REG <= 8'hb7;
        8'haa: OUT_REG <= 8'h62;
        8'hab: OUT_REG <= 8'h0e;
        8'hac: OUT_REG <= 8'haa;
        8'had: OUT_REG <= 8'h18;
        8'hae: OUT_REG <= 8'hbe;
        8'haf: OUT_REG <= 8'h1b;
        8'hb0: OUT_REG <= 8'hfc;
        8'hb1: OUT_REG <= 8'h56;
        8'hb2: OUT_REG <= 8'h3e;
        8'hb3: OUT_REG <= 8'h4b;
        8'hb4: OUT_REG <= 8'hc6;
        8'hb5: OUT_REG <= 8'hd2;
        8'hb6: OUT_REG <= 8'h79;
        8'hb7: OUT_REG <= 8'h20;
        8'hb8: OUT_REG <= 8'h9a;
        8'hb9: OUT_REG <= 8'hdb;
        8'hba: OUT_REG <= 8'hc0;
        8'hbb: OUT_REG <= 8'hfe;
        8'hbc: OUT_REG <= 8'h78;
        8'hbd: OUT_REG <= 8'hcd;
        8'hbe: OUT_REG <= 8'h5a;
        8'hbf: OUT_REG <= 8'hf4;
        8'hc0: OUT_REG <= 8'h1f;
        8'hc1: OUT_REG <= 8'hdd;
        8'hc2: OUT_REG <= 8'ha8;
        8'hc3: OUT_REG <= 8'h33;
        8'hc4: OUT_REG <= 8'h88;
        8'hc5: OUT_REG <= 8'h07;
        8'hc6: OUT_REG <= 8'hc7;
        8'hc7: OUT_REG <= 8'h31;
        8'hc8: OUT_REG <= 8'hb1;
        8'hc9: OUT_REG <= 8'h12;
        8'hca: OUT_REG <= 8'h10;
        8'hcb: OUT_REG <= 8'h59;
        8'hcc: OUT_REG <= 8'h27;
        8'hcd: OUT_REG <= 8'h80;
        8'hce: OUT_REG <= 8'hec;
        8'hcf: OUT_REG <= 8'h5f;
        8'hd0: OUT_REG <= 8'h60;
        8'hd1: OUT_REG <= 8'h51;
        8'hd2: OUT_REG <= 8'h7f;
        8'hd3: OUT_REG <= 8'ha9;
        8'hd4: OUT_REG <= 8'h19;
        8'hd5: OUT_REG <= 8'hb5;
        8'hd6: OUT_REG <= 8'h4a;
        8'hd7: OUT_REG <= 8'h0d;
        8'hd8: OUT_REG <= 8'h2d;
        8'hd9: OUT_REG <= 8'he5;
        8'hda: OUT_REG <= 8'h7a;
        8'hdb: OUT_REG <= 8'h9f;
        8'hdc: OUT_REG <= 8'h93;
        8'hdd: OUT_REG <= 8'hc9;
        8'hde: OUT_REG <= 8'h9c;
        8'hdf: OUT_REG <= 8'hef;
        8'he0: OUT_REG <= 8'ha0;
        8'he1: OUT_REG <= 8'he0;
        8'he2: OUT_REG <= 8'h3b;
        8'he3: OUT_REG <= 8'h4d;
        8'he4: OUT_REG <= 8'hae;
        8'he5: OUT_REG <= 8'h2a;
        8'he6: OUT_REG <= 8'hf5;
        8'he7: OUT_REG <= 8'hb0;
        8'he8: OUT_REG <= 8'hc8;
        8'he9: OUT_REG <= 8'heb;
        8'hea: OUT_REG <= 8'hbb;
        8'heb: OUT_REG <= 8'h3c;
        8'hec: OUT_REG <= 8'h83;
        8'hed: OUT_REG <= 8'h53;
        8'hee: OUT_REG <= 8'h99;
        8'hef: OUT_REG <= 8'h61;
        8'hf0: OUT_REG <= 8'h17;
        8'hf1: OUT_REG <= 8'h2b;
        8'hf2: OUT_REG <= 8'h04;
        8'hf3: OUT_REG <= 8'h7e;
        8'hf4: OUT_REG <= 8'hba;
        8'hf5: OUT_REG <= 8'h77;
        8'hf6: OUT_REG <= 8'hd6;
        8'hf7: OUT_REG <= 8'h26;
        8'hf8: OUT_REG <= 8'he1;
        8'hf9: OUT_REG <= 8'h69;
        8'hfa: OUT_REG <= 8'h14;
        8'hfb: OUT_REG <= 8'h63;
        8'hfc: OUT_REG <= 8'h55;
        8'hfd: OUT_REG <= 8'h21;
        8'hfe: OUT_REG <= 8'h0c;
        8'hff: OUT_REG <= 8'h7d;
      endcase
    end
  
    assign OUT_DATA = OUT_REG;
  
  endmodule
  